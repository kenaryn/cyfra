module main

import time
import util

fn main() {
    sw := time.new_stopwatch()

    get_stat()
}
